library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use work.opCodes_Pkg.ALL;

entity InstructionMemory is
    generic (
        N : integer := 8
    );
    port (
        addr       : in  STD_LOGIC_VECTOR(N-1 downto 0); 
        instr_out  : out STD_LOGIC_VECTOR(31 downto 0)  
    );
end InstructionMemory;

architecture Behavioral of InstructionMemory is

    signal instr_reg : STD_LOGIC_VECTOR(31 downto 0);
    -- Instruction memory array: each entry is a 32-bit instruction
    type instruction_mem_type is array(0 to 255) of STD_LOGIC_VECTOR(31 downto 0);
    signal instr_mem : instruction_mem_type := (
        
    0 => make_instr(OP_NOP, (others => '0'), (others => '0'), (others => '0')), --As a quick hacky fix, we need the first instruction to be nothing as it's skipped. 
    --------------------------------------------------
    --Here's where we can write our program
    -- the format of each instruction should be '[PC number] => marke_instr([OpCode], [arg1], [arg2], arg3]),' 
    -- If you want to refernce a register it needs to be in the form 'regcode_to_stdvec([register number])'
    -------------------------------------------------

    1 => make_instr(OP_MOV, x"01", (others => '0'), regcode_to_stdvec(R7)),
    2 => make_instr(OP_MOV, x"05", (others => '0'), regcode_to_stdvec(R0)),
    3 => make_instr(OP_MOV, x"00", (others => '0'), regcode_to_stdvec(R1)),
    4 => make_instr(OP_SUB, regcode_to_stdvec(R0), regcode_to_stdvec(R7), regcode_to_stdvec(R0)),
    5 => make_instr(OP_JGT, regcode_to_stdvec(R0), regcode_to_stdvec(R1), x"04"),
    6 => make_instr(OP_MOV, x"FF", (others => '0'), regcode_to_stdvec(R6)),




    --end program here
    -------------------------------------------------
        others => (others => '0') --All locations not defined in the program above will be zeroes.
    );

begin

    instr_out <= instr_mem(to_integer(unsigned(addr)));

end Behavioral;
